`timescale 1ns/1ps
import spi_config_pkg :: SPI_CLK_DIVIDE;
module spi_clk(
    input en,
    input logic sys_clk,
    output logic spi_clk
);



endmodule